
`define PACKET 10        // repeat in sequence


`define ADDR_WIDTH 32     
`define DATA_WIDTH 32
 
`define SEL 4
`define STR 4
